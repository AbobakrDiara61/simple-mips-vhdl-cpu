library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.ALL;

entity cpu is
 port(

 );
end cpu;

architecture behaviore of cpu is 
	-- signal section

	begin 
		process ()
		begin
		
		end process;
end behavioral

